class PySVObject;
chandle pysv_ptr;
endclass