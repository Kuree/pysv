import "DPI-C" function int simple_func(input int a,
                                        input int b,
                                        input int c);